entity MUXrf is
	port(
	ent1: in STD_LOGIC_VECTOR (4 downto 0);
	ent2: in STD_LOGIC_VECTOR (4 downto 0);
	sal_ out STD_LOGIC_VECTOR (4 downto 0)
	);
end MUXrf;

architecture MUXrf_arch of MUXrf is

end MUXrf_arch;