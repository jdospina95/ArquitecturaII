entity adderB is
	port(
	pcadd: in STD_LOGIC_VECTOR (31 downto 0);
	branchA: in STD_LOGIC_VECTOR (31 downto 0):
	resl: out STD_LOGIC_VECTOR (31 downto 0)
	);
end adderB

architecture adderB_arch of adderB is

end adderB_arch