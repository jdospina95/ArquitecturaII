entity instmemory is
	port(
	ent: in STD_LOGIC_VECTOR (31 downto 0);
	sal: in STD_LOGIC_VECTOR (31 downto 0));
end instmemory;

architecture instmemory_arch of instmemory is

end instmemory_arch